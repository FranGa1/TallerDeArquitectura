-------------------------------------------------------------------------------
--
-- Title       : pruebas
-- Design      : taller_de_arqui
-- Author      : franciscogaray
-- Company     : Facultad de Informatica UNLP
--
-------------------------------------------------------------------------------
--
-- File        : C:\My_Designs\taller_de_arqui\taller_de_arqui\src\pruebas.vhd
-- Generated   : Fri Sep 16 11:30:53 2022
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {pruebas} architecture {pruebas}}



entity pruebas is
end pruebas;

--}} End of automatically maintained section

architecture pruebas of pruebas is 
	signal c : integer;
begin

	 

end pruebas;
